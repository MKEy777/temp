`timescale 1ns / 1ps

/*
 * ģ��: SEE_Weight_BRAM
 * ����: 32-bit ��˫�˿� BRAM (1R1W)��
 * ְ��: �洢 SNN Ȩ�أ�֧�� 32-bit ���ȡ��
 */
module SEE_Weight_BRAM #(
    parameter DATA_W   = 32, 
    parameter ADDR_W   = 10, 
    parameter MEM_FILE = ""
)(
    input  wire                  clk,
    
    // �˿� A: ���˿� (-> SNN_Array_4PE)
    input  wire                  i_rd_en_a,
    input  wire [ADDR_W-1:0]     i_rd_addr_a,
    output reg signed [DATA_W-1:0] o_rd_data_a,

    // �˿� B: д�˿� (���ڼ���Ȩ��)
    input  wire                  i_wr_en_b,
    input  wire [ADDR_W-1:0]     i_wr_addr_b,
    input  wire signed [DATA_W-1:0] i_wr_data_b
);

    localparam MEM_DEPTH = 1 << ADDR_W;
    
    (* ram_style = "block" *) 
    reg [DATA_W-1:0] mem [0:MEM_DEPTH-1];

    initial begin
        if (MEM_FILE != "") begin
            $readmemh(MEM_FILE, mem);
        end
    end

    // �˿� A: ���߼� (ʱ��)
    always @(posedge clk) begin
        if (i_rd_en_a) begin
            o_rd_data_a <= mem[i_rd_addr_a];
        end
    end

    // �˿� B: д�߼� (ʱ��)
    always @(posedge clk) begin
        if (i_wr_en_b) begin
            mem[i_wr_addr_b] <= i_wr_data_b;
        end
    end

endmodule