`timescale 1ns / 1ps

/*
 * ģ��: PE_GALS_Wrapper [�ع���]
 * ����: GALS FSM, ʵ�� SNN �ĵ�λ�ۼӡ�
 * �ع�: �Ƴ��� o_bram_addr������� i_clk_en (ʱ��ʹ��)��
 */
module PE_GALS_Wrapper #(
    // Q1.7 Эͬ��Ʋ���
    parameter TIME_W   = 8,
    parameter WEIGHT_W = 8,
    
    // �ܹ�����
    parameter ADDR_W   = 10, // BRAM ��ַλ��
    parameter ACC_W    = 32  // 32-bit �ۼ��� (�����)
)(
    input  wire                 local_clk,
    input  wire                 rst_n,
    input  wire                 i_clk_en, // ** ����: ʱ��ʹ�� **

    // GALS �¼����� (�첽����)
    input  wire                 i_aer_req,
    input  wire signed [TIME_W-1:0] i_aer_time, // 8-bit (t_i)
    input  wire [ADDR_W-1:0]        i_aer_addr,
    
    // SNN FSM ���Ʋ���
    input  wire signed [TIME_W-1:0] i_t_min,    // 8-bit (t_min)
    input  wire                 i_reset_potential,

    // GALS ������� (-> Collector)
    output reg                  o_done_req,
    input  wire                 i_done_ack,

    // ר�� BRAM �ӿ�
    output reg                  o_bram_en,
    // [���Ƴ�] o_bram_addr �˿�
    input  wire signed [WEIGHT_W-1:0] i_bram_data, // 8-bit (W_ij)

    // ��λ��� (-> SNN_Engine)
    output wire signed [ACC_W-1:0]  o_potential_j // 32-bit (V_j)
);

    // GALS FSM ״̬����
    localparam S_IDLE       = 4'b0000;
    localparam S_LATCH_AER  = 4'b0001; // C1: ����, �ύBRAM En
    localparam S_READ_BRAM  = 4'b0010; // C2: ��BRAM, ���� (t_i - t_min)
    localparam S_COMPUTE    = 4'b0011; // C3: BRAM������Ч, ���� (t_diff * W_ij)
    localparam S_ACCUMULATE = 4'b0100; // C4: �ۼ�, ���� o_done_req
    localparam S_WAIT_ACK   = 4'b0101; // C5: �ȴ� Collector ȷ��

    reg [3:0] state, next_state;

    // �ڲ�����·���Ĵ���
    reg signed [ACC_W-1:0]   V_j_reg;
    reg signed [TIME_W-1:0]  latched_aer_time;
    // [���Ƴ�] latched_aer_addr
    
    // ��ˮ�߽׶μĴ���
    reg signed [TIME_W:0]    p2_time_diff;   // (t_i - t_min) -> 9b
    reg signed [ACC_W-1:0]   p3_mult_result; // (t_diff * W_ij) -> 17b (��չ)
    
    assign o_potential_j = V_j_reg;

    // 1. FSM ״̬�� (����߼�)
    // (�ⲿ�ֲ���Ҫʱ��ʹ�ܣ����ֲ���)
    always @(*) begin
        next_state  = state;
        o_done_req  = 1'b0;
        o_bram_en   = 1'b0;

        case (state)
            S_IDLE: begin
                if (i_aer_req)
                    next_state = S_LATCH_AER;
            end
            
            S_LATCH_AER: begin
                o_bram_en = 1'b1; // C1: ���ύ BRAM ��ʹ��
                next_state = S_READ_BRAM;
            end

            S_READ_BRAM: begin
                next_state = S_COMPUTE;
            end

            S_COMPUTE: begin
                next_state = S_ACCUMULATE;
            end
            
            S_ACCUMULATE: begin
                o_done_req = 1'b1;
                next_state = S_WAIT_ACK;
            end
            
            S_WAIT_ACK: begin
                o_done_req = 1'b1;
                if (i_done_ack)
                    next_state = S_IDLE;
            end

            default: begin
                next_state = S_IDLE;
            end
        endcase
    end

    // 2. FSM ������·�� (ʱ���߼�)
    // ** �ؼ�: ����ʱ���߼��������� i_clk_en ���� **
    always @(posedge local_clk or negedge rst_n) begin
        if (!rst_n) begin
            state            <= S_IDLE;
            V_j_reg          <= {ACC_W{1'b0}};
            latched_aer_time <= {TIME_W{1'b0}};
            p2_time_diff     <= 0;
            p3_mult_result   <= 0;
        end 
        // ** ֻ���� rst_n ��Ч�� i_clk_en ��Чʱ����ִ��ʱ���߼� **
        else if (i_clk_en) begin 
            
            state <= next_state;
            
            if (i_reset_potential) begin
                V_j_reg <= {ACC_W{1'b0}};
            end

            // ����·����ˮ��
            case (state)
                S_LATCH_AER: begin 
                    // C1: ����ʱ�� (������Ҫ�����ַ)
                    latched_aer_time <= i_aer_time;
                end

                S_READ_BRAM: begin 
                    // C2: ���� (t_i - t_min)
                    p2_time_diff <= $signed(latched_aer_time) - $signed(i_t_min);
                end
                
                S_COMPUTE: begin 
                    // C3: ���� (t_diff * W_ij)
                    p3_mult_result <= $signed(p2_time_diff) * $signed(i_bram_data);
                end
                
                S_ACCUMULATE: begin 
                    // C4: �ۼ� (V_j_reg += product)
                    if (!i_reset_potential)
                        V_j_reg <= V_j_reg + p3_mult_result;
                end
            endcase
        end
    end

endmodule