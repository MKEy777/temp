`timescale 1ns / 1ps

module ram_sync #(
    parameter DATA_WIDTH = 24,
    parameter ADDR_WIDTH = 10,
    parameter MEM_FILE   = ""    
)(
    input  wire                  clk,
    
    // д�˿� (Port A)
    input  wire                  wr_en,
    input  wire [ADDR_WIDTH-1:0] wr_addr,
    input  wire [DATA_WIDTH-1:0] wr_data,
    
    // ���˿� (Port B)
    input  wire                  rd_en,
    input  wire [ADDR_WIDTH-1:0] rd_addr,
    output reg  [DATA_WIDTH-1:0] rd_data
);

    localparam MEM_DEPTH = 1 << ADDR_WIDTH;

    // ǿ���ƶ�Ϊ Block RAM
    (* ram_style = "block" *) 
    reg [DATA_WIDTH-1:0] mem [0:MEM_DEPTH-1];

    // ��ʼ�� (ͨ�����ڷ��棬FPGA�ϵ��ʼֵ)
    integer i;
    initial begin
        if (MEM_FILE != "") begin
            $readmemh(MEM_FILE, mem);
        end else begin
            // ���û���ļ�����ʼ��Ϊȫ0 (����SNNĤ��λ����Ҫ)
            for (i = 0; i < MEM_DEPTH; i = i + 1) begin
                mem[i] = 0;
            end
        end
    end

    // д�߼� (Port A)
    always @(posedge clk) begin
        if (wr_en) begin
            mem[wr_addr] <= wr_data;
        end
    end

    // ���߼� (Port B)
    always @(posedge clk) begin
        if (rd_en) begin
            rd_data <= mem[rd_addr];
        end
    end

endmodule