`timescale 1ns / 1ps

/*
 * ģ��: GALS_Encoder_Unit
 * ����: GALS �Ž������� ANN ����ֵ (Q1.7) ת��Ϊ SNN ����ʱ�� (Q1.7)��
 * �㷨: t_i = T_MAX - ((x - K_MIN) >> K_SHIFT)
 */
module GALS_Encoder_Unit #(
    // �ܹ�����
    parameter VEC_LEN       = 160, // SNN ����ά�� (8x4x5)
    parameter PIXEL_VEC_LEN = 8,   // ANN �ں� FSM ÿ�η��͵�ͨ����
    parameter NUM_PIXELS    = 20,  // VEC_LEN / PIXEL_VEC_LEN
    parameter DATA_W        = 8,   // Q1.7 ����ֵ (���� ANN)
    parameter TIME_W        = 8,   // Q1.7 ����ʱ�� (���� SNN)
    
    // Q1.7 ���볣�� (�������ѵ��)
    parameter signed [DATA_W-1:0] T_MAX_Q17 = 127,
    parameter signed [DATA_W-1:0] K_MIN_Q17 = -128,
    parameter SHIFT_BITS    = 2    // ʾ��ֵ
)(
    input  wire                      local_clk,
    input  wire                      rst_n,

    // GALS ���� (���� ULG_Coordinator)
    input  wire                      i_data_req,
    output reg                       o_data_ack,
    input  wire signed [PIXEL_VEC_LEN*DATA_W-1:0] i_data_bus, 

    // AER �㲥���� (-> SNN_Engine)
    output reg                       o_aer_req,
    input  wire                      i_aer_ack,
    output reg signed [TIME_W-1:0]   o_aer_time,
    output reg [$clog2(VEC_LEN)-1:0] o_aer_addr,
    
    output wire                      o_busy,
    output wire                      o_encoder_done
);

    // FSM ״̬
    localparam S_IDLE       = 3'b000;
    localparam S_CALC_LOAD  = 3'b001; 
    localparam S_SEND_SPIKE = 3'b010;
    localparam S_FINISHING  = 3'b011;
    reg [2:0] state, next_state;

    // ������
    reg [$clog2(NUM_PIXELS)-1:0]    pixel_receive_cnt; // 0-19
    reg [$clog2(PIXEL_VEC_LEN)-1:0] channel_send_cnt;  // 0-7
    
    // �ڲ��Ĵ���
    reg signed [TIME_W-1:0] current_pixel_spikes [0:PIXEL_VEC_LEN-1];
    wire signed [TIME_W-1:0] calculated_spikes [0:PIXEL_VEC_LEN-1];

    // Q1.7 �����㷨 (����߼�)
    genvar i;
    generate
        for (i = 0; i < PIXEL_VEC_LEN; i = i + 1) begin : PIXEL_ENCODE_LOGIC
            wire signed [DATA_W-1:0] x_q;
            wire signed [DATA_W:0]   x_sub;     // (x - K_MIN) -> 9b
            wire signed [DATA_W:0]   x_shift;   // (x_sub >> K_SHIFT)
            wire signed [DATA_W-1:0] x_clamped; // clamp(x_shift, 0, 127)
            
            assign x_q = i_data_bus[(i+1)*DATA_W-1 -: DATA_W];
            
            // �㷨 1: (x - K_MIN_Q17)
            assign x_sub = $signed(x_q) - $signed(K_MIN_Q17);
            
            // �㷨 2: (x_sub >>> K_SHIFT) (��������)
            assign x_shift = x_sub >>> SHIFT_BITS;
            
            // �㷨 3: clamp(..., 0, T_MAX_Q17)
            assign x_clamped = (x_shift < 0) ? 0 : 
                               (x_shift > T_MAX_Q17) ? T_MAX_Q17 : 
                               x_shift[DATA_W-1:0];
                               
            // �㷨 4: t_i = T_MAX - clamped_norm_x
            assign calculated_spikes[i] = T_MAX_Q17 - x_clamped;
        end
    endgenerate

    // 1. FSM (����߼�)
    always @(*) begin
        next_state = state;
        o_aer_req  = 1'b0;
        o_aer_time = {TIME_W{1'bx}};
        o_aer_addr = {$clog2(VEC_LEN){1'bx}};
        o_data_ack = 1'b0;

        case (state)
            S_IDLE: begin
                if (i_data_req) begin
                    o_data_ack = 1'b1;
                    next_state = S_CALC_LOAD;
                end
            end
            
            S_CALC_LOAD: begin
                o_data_ack = 1'b1;
                if (!i_data_req)
                    next_state = S_SEND_SPIKE;
            end

            S_SEND_SPIKE: begin
                // ��������Ƿ���Ч (������Ч����)
                if (current_pixel_spikes[channel_send_cnt] < T_MAX_Q17) begin
                    o_aer_req  = 1'b1;
                    o_aer_time = current_pixel_spikes[channel_send_cnt];
                    o_aer_addr = (pixel_receive_cnt * PIXEL_VEC_LEN) + channel_send_cnt;
                    
                    if (i_aer_ack) begin // ���ֳɹ�, ׼����һ��
                        if (channel_send_cnt == PIXEL_VEC_LEN - 1)
                            next_state = (pixel_receive_cnt == NUM_PIXELS - 1) ?
                                         S_FINISHING : S_IDLE;
                        else
                            next_state = S_SEND_SPIKE;
                    end else
                        next_state = S_SEND_SPIKE; // ���� req, �ȴ� ack
                end else begin
                    // ������Ч���� (>= T_MAX_Q17)
                    if (channel_send_cnt == PIXEL_VEC_LEN - 1)
                        next_state = (pixel_receive_cnt == NUM_PIXELS - 1) ?
                                     S_FINISHING : S_IDLE;
                    else
                        next_state = S_SEND_SPIKE;
                end
            end

            S_FINISHING: next_state = S_IDLE;
            default:     next_state = S_IDLE;
        endcase
    end
    
    // 2. FSM (ʱ���߼�)
    integer ch;
    always @(posedge local_clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_IDLE;
            pixel_receive_cnt <= 0;
            channel_send_cnt <= 0;
            for (ch = 0; ch < PIXEL_VEC_LEN; ch = ch + 1)
                current_pixel_spikes[ch] <= T_MAX_Q17; // ��λΪ "��Ч"
        end else begin
            state <= next_state;

            case (state)
                S_IDLE: begin
                    if (next_state == S_CALC_LOAD) begin
                        if (pixel_receive_cnt == NUM_PIXELS - 1)
                            pixel_receive_cnt <= 0;
                        else
                            pixel_receive_cnt <= pixel_receive_cnt + 1;
                    end
                end

                S_CALC_LOAD: begin
                    if (next_state == S_SEND_SPIKE) begin
                        for (ch = 0; ch < PIXEL_VEC_LEN; ch = ch + 1)
                            current_pixel_spikes[ch] <= calculated_spikes[ch];
                        channel_send_cnt <= 0;
                    end
                end
                
                S_SEND_SPIKE: begin
                    // ���� (���屻����) �� (���巢�ͳɹ�) ʱ���ŵ���������
                    if (current_pixel_spikes[channel_send_cnt] >= T_MAX_Q17 || (o_aer_req && i_aer_ack)) begin
                        if (channel_send_cnt != PIXEL_VEC_LEN - 1)
                            channel_send_cnt <= channel_send_cnt + 1;
                    end
                end
                
                S_FINISHING: begin
                    pixel_receive_cnt <= 0;
                    channel_send_cnt  <= 0;
                end
            endcase
        end
    end
    
    assign o_busy = (state != S_IDLE);
    assign o_encoder_done = (state == S_FINISHING); 

endmodule