`timescale 1ns/1ps
`default_nettype wire

// MACƫ�ô���Ԫģ��
// ���ܣ����ƫ�üӷ���������ս��
module mac_bias_unit #(
    parameter DATA_WIDTH = 16,    // MAC�������λ��
    parameter BIAS_WIDTH = 16,    // ƫ��λ��
    parameter OUT_WIDTH = 18      // ���λ�����Ǽӷ������
)(
    input  wire                    clk,           // ʱ��
    input  wire                    rst_n,         // ��λ������Ч
    input  wire                    valid_in,      // ������Ч�ź�
    input  wire [DATA_WIDTH-1:0]   mac_data,      // MAC�������
    input  wire [BIAS_WIDTH-1:0]   bias_data,     // ƫ������
    output wire [OUT_WIDTH-1:0]    result_data,   // ���ս��
    output wire                    valid_out      // �����Ч�ź�
);

// �ڲ��źŶ���
wire signed [OUT_WIDTH-1:0] bias_add_result;

// ƫ�üӷ�
// ʹ�� $signed() ��ʽ��֪�ۺ��������з��żӷ�
assign bias_add_result = $signed(mac_data) + $signed(bias_data);

// ��ˮ�߼Ĵ����ź�
reg [OUT_WIDTH-1:0] result_data_reg;
reg                 valid_out_reg;

// ��ʱ���߼� - ������ˮ��
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        result_data_reg <= 0;
        valid_out_reg <= 0;
    end else begin
        result_data_reg <= bias_add_result;
        valid_out_reg <= valid_in;
    end
end

// �������
assign result_data = result_data_reg;
assign valid_out = valid_out_reg;

endmodule