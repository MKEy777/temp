`timescale 1ns / 1ps

/*
 * ģ��: Feature_Map_Buffer_1W3R
 * ����: 1д3�� (1W3R) ͬ��RAM��
 * ʵ��: ͨ�����ݸ��� (Replication) ʵ�֡�
 * C1 FSM ������3���ڲ�RAMд�룬P1/P2/P3 ���Զ�ȡ1����
 */
module Feature_Map_Buffer_1W3R #(
    parameter DATA_WIDTH = 8,
    parameter ADDR_WIDTH = 10,
    parameter RAM_DEPTH  = 1 << ADDR_WIDTH
)(
    input  wire                      clk,

    // --- �˿� A: д�˿� (���� C1 FSM) ---
    input  wire                      i_wr_en,
    input  wire [ADDR_WIDTH-1:0]     i_wr_addr,
    input  wire signed [DATA_WIDTH-1:0]  i_wr_data,

    // --- �˿� A: ���˿� (���� P1: Main Path) ---
    input  wire                      i_rd_en_a,
    input  wire [ADDR_WIDTH-1:0]     i_rd_addr_a,
    output reg signed [DATA_WIDTH-1:0]  o_rd_data_a,

    // --- �˿� B: ���˿� (���� P2: Channel Gate) ---
    input  wire                      i_rd_en_b,
    input  wire [ADDR_WIDTH-1:0]     i_rd_addr_b,
    output reg signed [DATA_WIDTH-1:0]  o_rd_data_b,

    // --- �˿� C: ���˿� (���� P3: Spatial Gate) ---
    input  wire                      i_rd_en_c,
    input  wire [ADDR_WIDTH-1:0]     i_rd_addr_c,
    output reg signed [DATA_WIDTH-1:0]  o_rd_data_c
);

    // ʵ���� 3 �������� BRAM
    (* ram_style = "block" *)
    reg [DATA_WIDTH-1:0] mem_a [0:RAM_DEPTH-1];
    
    (* ram_style = "block" *)
    reg [DATA_WIDTH-1:0] mem_b [0:RAM_DEPTH-1];
    
    (* ram_style = "block" *)
    reg [DATA_WIDTH-1:0] mem_c [0:RAM_DEPTH-1];

    // --- �˿� A: д�߼� (ͬʱд������ BRAM) ---
    always @(posedge clk) begin
        if (i_wr_en) begin
            mem_a[i_wr_addr] <= i_wr_data;
            mem_b[i_wr_addr] <= i_wr_data;
            mem_c[i_wr_addr] <= i_wr_data;
        end
    end

    // --- �˿� A, B, C: ���߼� (���Զ�ȡ) ---
    always @(posedge clk) begin
        if (i_rd_en_a) begin
            o_rd_data_a <= mem_a[i_rd_addr_a];
        end
        
        if (i_rd_en_b) begin
            o_rd_data_b <= mem_b[i_rd_addr_b];
        end
        
        if (i_rd_en_c) begin
            o_rd_data_c <= mem_c[i_rd_addr_c];
        end
    end

endmodule