`timescale 1ns / 1ps

/*
 * ģ��: GALS_Accelerator_Top
 * ����: GALS���ANN-SNN�������Ķ����װ��
 * ְ��:
 * 1. ���� ANN_Engine, GALS_Encoder_Unit, SNN_Engine��
 * 2. ���Ӷ��� GALS �첽���ֽӿڡ�
 * 3. ��������Ӳ��������
 * 4. ��¶���ݺ�Ȩ��/ƫ�õĶ��� I/O��
 */
module GALS_Accelerator_Top #(
    // --- ���� Q1.7 ���� ---
    parameter DATA_W    = 8,   // ����/Ȩ�� (Q1.7)
    parameter TIME_W    = 8,   // ����ʱ�� (Q1.7)
    parameter WEIGHT_W  = 8,   // SNN Ȩ�� (Q1.7)
    parameter ACC_W     = 32,  // 32-bit �ۼ���
    
    // --- ������� ---
    parameter K_DIM     = 3,   // 3x3 �����
    
    // --- ANN C1 ���� (���� QAT.py) ---
    parameter C1_IN_CH  = 4,
    parameter C1_OUT_CH = 8,
    parameter C1_IMG_W  = 9,
    parameter C1_IMG_H  = 8,
    
    // --- ANN C2 ���� (���� QAT.py) ---
    parameter C2_IN_CH  = 8,   // C1_OUT_CH
    parameter C2_IMG_W  = 5,   // C1 ���/������Ľ��
    parameter C2_IMG_H  = 4,
    
    // --- ANN Requantize ���� ---
    parameter C1_BIAS_W     = 32,
    parameter C1_SHIFT_BITS = 14, // ʾ��
    
    // --- SNN ���� (���� QAT.py �� SNN_Engine.v) ---
    parameter SNN_IN_LEN     = 160, // 8 (C2_IN_CH) * 5 * 4 = 160
    parameter DENSE1_NEURONS = 64,
    parameter DENSE2_NEURONS = 32,
    parameter DENSE3_NEURONS = 3,
    parameter NUM_ARRAYS     = 16,  // 64 PE / 4 PE-per-Array
    
    // --- ��ַ���߿�� ---
    parameter FM_ADDR_W = 10,  // ����ͼ BRAM ��ַ
    parameter ADDR_W    = 10   // SNN BRAM ��ַ
)(
    input  wire                      clk,
    input  wire                      rst_n,

    // --- ANN ��������ӿ� ---
    input  wire                      i_data_req,    // ��������һ֡ (�����ⲿ)
    input  wire signed [C1_IN_CH*DATA_W-1:0] i_data_flat, // ANN ����������
    output wire                      o_data_ack,    // ȷ���յ�ANN����

    // --- SNN ������ƽӿ� ---
    input  wire                      i_accelerator_start, // ���� SNN (�����ⲿ)
    output wire                      o_accelerator_done,  // SNN ���
    output wire [$clog2(DENSE3_NEURONS)-1:0] o_predicted_class, // SNN ���

    // --- Ȩ��/ƫ�� ROM �ӿ� (�����ⲿ) ---
    
    // ANN C1 (DSC)
    input  wire signed [C1_IN_CH*K_DIM*K_DIM*DATA_W-1:0] i_kernel_c1_dw,
    input  wire signed [C1_OUT_CH*C1_IN_CH*DATA_W-1:0] i_kernel_c1_pw,
    input  wire signed [C1_BIAS_W-1:0]                 i_bias_c1_requant_dw,
    input  wire signed [C1_BIAS_W-1:0]                 i_bias_c1_requant_pw,
    
    // ANN C2 (ULG)
    input  wire signed [C2_IN_CH*K_DIM*K_DIM*DATA_W-1:0] i_kernel_c2_p1,
    input  wire signed [C2_IN_CH*C2_IN_CH*DATA_W-1:0] i_kernel_c2_p2,
    input  wire signed [K_DIM*K_DIM*DATA_W-1:0] i_kernel_c2_p3,
    
    // SNN �����ֵ (�����ⲿ ROM)
    /*
     * ע: SNN_Engine ���� i_snn_threshold_data �˿�����ȷ��ʱ��
     * (�� SNN_Engine �ڲ��� Intermediate_Buffer_Encoder ����) 
     * Я����ȷ����ֵ D_i��
     * ��ʵ��ϵͳ�У�����Ҫһ�� ROM�����ַ�� SNN_Engine ��
     * �ڲ��ź����� (�õ�ַ�˿��� SNN_Engine.v ��δ������)��
     * �˴����ǽ���¶ SNN_Engine.v ��������ݶ˿ڡ�
     */
    input  wire signed [WEIGHT_W-1:0] i_snn_threshold_data
);

    // =========================================================================
    // 1. GALS ��������
    // =========================================================================
    
    // --- �ӿ� 1: ANN_Engine -> GALS_Encoder_Unit ---
    // (ANN ���� Q1.7 ������)
    wire        ann_to_enc_req;
    wire        ann_to_enc_ack;
    wire signed [C2_IN_CH*DATA_W-1:0] ann_to_enc_data; // (8-channel wide)
    
    // --- �ӿ� 2: GALS_Encoder_Unit -> SNN_Engine ---
    // (Encoder �㲥 Q1.7 AER ����)
    wire        enc_to_snn_req;
    wire        enc_to_snn_ack;
    wire        enc_to_snn_done;
    wire signed [TIME_W-1:0] enc_to_snn_time;
    
    // ��ַ����ƥ��
    localparam SNN_ADDR_W = $clog2(SNN_IN_LEN); // 8-bit (for 160)
    wire [SNN_ADDR_W-1:0] enc_to_snn_addr_raw;
    wire [ADDR_W-1:0]     enc_to_snn_addr_padded;
    
    // SNN_Engine ���� [ADDR_W-1:0] ����, 
    // GALS_Encoder ��� [$clog2(VEC_LEN)-1:0]
    assign enc_to_snn_addr_padded = { {(ADDR_W - SNN_ADDR_W){1'b0}}, enc_to_snn_addr_raw };


    // =========================================================================
    // 2. ���� GALS ģ��
    // =========================================================================

    // --- ģ�� 1: ANN ǰ������ ---
    ANN_Engine #(
        .DATA_W    ( DATA_W    ), .ACC_W     ( ACC_W     ), .K_DIM     ( K_DIM     ),
        .C1_IN_CH  ( C1_IN_CH  ), .C1_OUT_CH ( C1_OUT_CH ), .C1_IMG_W  ( C1_IMG_W  ),
        .C1_IMG_H  ( C1_IMG_H  ), .C2_IN_CH  ( C2_IN_CH  ), .C2_IMG_W  ( C2_IMG_W  ),
        .C2_IMG_H  ( C2_IMG_H  ), .FM_ADDR_W ( FM_ADDR_W ), .C1_BIAS_W ( C1_BIAS_W ),
        .C1_SHIFT_BITS( C1_SHIFT_BITS )
    ) ann_engine_inst (
        .clk        ( clk ),
        .rst_n      ( rst_n ),
        
        .i_data_req ( i_data_req ),
        .i_data_flat( i_data_flat ),
        .o_data_ack ( o_data_ack ),

        .o_encoder_req     ( ann_to_enc_req ),
        .i_encoder_ack     ( ann_to_enc_ack ),
        .o_encoder_data_flat( ann_to_enc_data ),
        
        .i_kernel_c1_dw      ( i_kernel_c1_dw ),
        .i_kernel_c1_pw      ( i_kernel_c1_pw ),
        .i_bias_c1_requant_dw( i_bias_c1_requant_dw ),
        .i_bias_c1_requant_pw( i_bias_c1_requant_pw ),
        .i_kernel_c2_p1      ( i_kernel_c2_p1 ),
        .i_kernel_c2_p2      ( i_kernel_c2_p2 ),
        .i_kernel_c2_p3      ( i_kernel_c2_p3 )
    );

    // --- ģ�� 2: GALS �Ž��� (ANN -> SNN) ---
  
    localparam ENCODER_PIXEL_VEC_LEN = C2_IN_CH;
    localparam ENCODER_NUM_PIXELS    = SNN_IN_LEN / ENCODER_PIXEL_VEC_LEN;
    
    GALS_Encoder_Unit #(
        .VEC_LEN       ( SNN_IN_LEN ),
        .PIXEL_VEC_LEN ( ENCODER_PIXEL_VEC_LEN ),
        .NUM_PIXELS    ( ENCODER_NUM_PIXELS ),
        .DATA_W        ( DATA_W ),
        .TIME_W        ( TIME_W ),
        

        .T_MAX_Q17 ( 8'd127 ),
        .K_MIN_Q17 ( -8'd128 ),
        .SHIFT_BITS( 2 )
    ) gals_encoder_inst (
        .local_clk ( clk ),
        .rst_n     ( rst_n ),

        // ���� ANN_Engine
        .i_data_req( ann_to_enc_req ),
        .o_data_ack( ann_to_enc_ack ),
        .i_data_bus( ann_to_enc_data ), 

        // ���� SNN_Engine
        .o_aer_req     ( enc_to_snn_req ),
        .i_aer_ack     ( enc_to_snn_ack ),
        .o_aer_time    ( enc_to_snn_time ),
        .o_aer_addr    ( enc_to_snn_addr_raw ),
        .o_encoder_done( enc_to_snn_done ),
        
        .o_busy ( /* δ���� */ )
    );

    // --- ģ�� 3: SNN ������� ---
    SNN_Engine #(
        .TIME_W      ( TIME_W ),
        .WEIGHT_W    ( WEIGHT_W ),
        .ACC_W       ( ACC_W ),
        .ADDR_W      ( ADDR_W ),
        .NUM_ARRAYS  ( NUM_ARRAYS ),
        .SNN_IN_LEN  ( SNN_IN_LEN ),
        .DENSE1_NEURONS ( DENSE1_NEURONS ),
        .DENSE2_NEURONS ( DENSE2_NEURONS ),
        .DENSE3_NEURONS ( DENSE3_NEURONS ),
        
        // BRAM ƫ���� (���� SNN_Engine.v Ĭ��ֵ)
        .BRAM_OFFSET_D1 ( 10'd0 ),
        .BRAM_OFFSET_D2 ( 10'd160 ), // SNN_IN_LEN
        .BRAM_OFFSET_D3 ( 10'd224 ), // 160 + 64
        
        // t_min (���� SNN_Engine.v Ĭ��ֵ)
        .T_MIN_D1_Q17 ( 8'd0 ),
        .T_MIN_D2_Q17 ( 8'd20 ),
        .T_MIN_D3_Q17 ( 8'd40 )
    ) snn_engine_inst (
        .local_clk ( clk ),
        .rst_n     ( rst_n ),

        // �������
        .i_accelerator_start( i_accelerator_start ),
        .o_accelerator_done ( o_accelerator_done ),
        .o_predicted_class  ( o_predicted_class ),

        // ���� GALS_Encoder_Unit
        .i_enc_aer_req    ( enc_to_snn_req ),
        .i_enc_aer_time   ( enc_to_snn_time ),
        .i_enc_aer_addr   ( enc_to_snn_addr_padded ), // ʹ������ĵ�ַ
        .i_enc_done       ( enc_to_snn_done ),
        .o_enc_aer_ack    ( enc_to_snn_ack ),

        // ��ֵ ROM �ӿ�
        .i_threshold_data ( i_snn_threshold_data )
    );

endmodule