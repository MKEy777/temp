`timescale 1ns / 1ps

/*
 * ģ��: arithmetic_unit
 * ����: ͬ����ˮ�߳˷��� (Q1.7 * Q1.7 => Q1.7)
 * ��Ϊ: 1. (Stage 1) A * B
 * 2. (Stage 2) (A*B) >>> 7 (�ض���) + ����
 * ����: ULG_Coordinator (C2) ʵ�� (A*B)*C �ں�
 */
module arithmetic_unit #(
    parameter DATA_W     = 8,   // int8 (Q1.7)
    parameter MULT_W     = 16,  // DATA_W * 2
    parameter SHIFT_BITS = 7    // Q2.14 -> Q1.7 (14-7=7)
) (
    input wire                      clk,
    input wire                      rst_n,
    input wire                      i_valid,
    input wire signed [DATA_W-1:0]  i_data_a,
    input wire signed [DATA_W-1:0]  i_data_b,
    
    output reg signed [DATA_W-1:0] o_data,
    output reg                      o_valid
);

    // int8 ���ͷ�Χ
    localparam Q_MIN = -(2**(DATA_W-1));      // -128
    localparam Q_MAX = (2**(DATA_W-1)) - 1;  //  127

    // --- ��ˮ�߼Ĵ������� ---

    // Pipeline Stage 1: �˷����
    reg p1_valid;
    reg signed [MULT_W-1:0] p1_mult_result; // 8b * 8b = 16b

    // Stage 2: ����߼�
    wire signed [MULT_W-1:0] shifted_result;
    
    // Q2.14 (16b) -> Qx.7 (16b)
    assign shifted_result = p1_mult_result >>> SHIFT_BITS;


    // --- ��ˮ���߼� ---

    // Stage 1: �˷�
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            p1_valid       <= 1'b0;
            p1_mult_result <= {MULT_W{1'b0}};
        end else begin
            p1_valid <= i_valid;
            if (i_valid) begin
                // ʹ�� DSP ��Դִ���з��ų˷�
                p1_mult_result <= $signed(i_data_a) * $signed(i_data_b);
            end
        end
    end

    // Stage 2: �ض���(��λ) �� ����
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            o_valid <= 1'b0;
            o_data  <= {DATA_W{1'b0}};
        end else begin
            o_valid <= p1_valid;
            
            if (p1_valid) begin
                // 1. ���ͼ�� (Saturation)
                if (shifted_result < Q_MIN) begin
                    o_data <= Q_MIN;
                end else if (shifted_result > Q_MAX) begin
                    o_data <= Q_MAX;
                // 2. ��ֵ
                end else begin
                    // ��ȡ��8λ (Qx.7 -> Q1.7)
                    o_data <= shifted_result[DATA_W-1:0];
                end
            end else begin
                o_data <= {DATA_W{1'b0}};
            end
        end
    end

endmodule