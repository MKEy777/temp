`timescale 1ns / 1ps

/*
 * ģ��: PE_GALS_Wrapper (SNN ����Ԫ)
 * ����: GALS FSM��ʵ��SNN��O(1)�¼�����
 * ��Ϊ:
 * 1. �첽���� (i_aer_req)
 * 2. ����AER���� (i_aer_addr, i_aer_time)
 * 3. ͬ���� BRAM (o_bram_addr <- i_aer_addr)
 * 4. ͬ������ (V_j_reg <= V_j_reg + (i_aer_time * W[i,j]))
 * 5. �첽���� (o_done_req -> i_done_ack)
 */
module PE_GALS_Wrapper #(
    parameter TIME_W   = 32, // ����ʱ��λ�� (���� GALS_Encoder)
    parameter WEIGHT_W = 8,  // Ȩ��λ�� (int8)
    parameter ADDR_W   = 9,  // BRAM ��ַλ�� (e.g., clog2(320))
    parameter ACC_W    = 48  // �ۼ���λ�� (ƥ�� ArgMax_Unit)
)(
    input  wire                      local_clk,
    input  wire                      rst_n,

    // --- ȫ���첽�¼����� (���� Encoder) ---
    input  wire                      i_aer_req,
    input  wire signed [TIME_W-1:0]  i_aer_time,
    input  wire [ADDR_W-1:0]         i_aer_addr,
    
    // --- PE������� (-> Collector) ---
    output reg                       o_done_req,
    input  wire                      i_done_ack,

    // --- ר�� BRAM �ӿ� (-> SEE_Weight_BRAM_j) ---
    output reg                       o_bram_en,
    output reg [ADDR_W-1:0]          o_bram_addr,
    input  wire signed [WEIGHT_W-1:0] i_bram_data, // W[i, j]

    // --- ��λ��λ����� (-> SNN_Engine / ArgMax_Unit) ---
    input  wire                      i_reset_potential, // ��SNN_Engine����
    output wire signed [ACC_W-1:0]   o_potential_j
);

    // --- FSM ״̬���� ---
    localparam S_IDLE       = 3'b000;
    localparam S_LATCH_AER  = 3'b001;
    localparam S_READ_BRAM  = 3'b010;
    localparam S_COMPUTE    = 3'b011;
    localparam S_SEND_DONE  = 3'b100;
    localparam S_WAIT_ACK   = 3'b101;

    reg [2:0] state, next_state;

    // --- �ڲ��Ĵ��� ---
    reg signed [ACC_W-1:0]   V_j_reg;
    reg signed [TIME_W-1:0]  latched_aer_time;
    reg [ADDR_W-1:0]         latched_aer_addr;
    reg signed [ACC_W-1:0]   mult_result;
    
    assign o_potential_j = V_j_reg;

    // --- ״̬�� (����߼�) ---
    always @(*) begin
        next_state  = state;
        o_done_req  = 1'b0;
        o_bram_en   = 1'b0;
        o_bram_addr = latched_aer_addr;
        
        case (state)
            S_IDLE: begin
                if (i_aer_req) begin
                    next_state = S_LATCH_AER;
                end
            end
            
            S_LATCH_AER: begin
                // ������������
                next_state = S_READ_BRAM;
            end

            S_READ_BRAM: begin
                // ���� BRAM ��
                o_bram_en = 1'b1;
                next_state = S_COMPUTE;
            end

            S_COMPUTE: begin
                // BRAM ���� (W[i,j]) �ڴ�ʱ��������Ч
                // ���㹱�ײ��ۼ�
                next_state = S_SEND_DONE;
            end
            
            S_SEND_DONE: begin
                o_done_req = 1'b1;
                next_state = S_WAIT_ACK;
            end
            
            S_WAIT_ACK: begin
                o_done_req = 1'b1;
                if (i_done_ack) begin
                    next_state = S_IDLE;
                end
            end

            default: begin
                next_state = S_IDLE;
            end
        endcase
    end

    // --- ״̬��������·�� (ʱ���߼�) ---
    always @(posedge local_clk or negedge rst_n) begin
        if (!rst_n) begin
            state            <= S_IDLE;
            V_j_reg          <= {ACC_W{1'b0}};
            latched_aer_time <= {TIME_W{1'b0}};
            latched_aer_addr <= {ADDR_W{1'b0}};
            mult_result      <= {ACC_W{1'b0}};
        end else begin
            state <= next_state;

            if (i_reset_potential) begin
                V_j_reg <= {ACC_W{1'b0}};
            end

            case (state)
                S_LATCH_AER: begin
                    latched_aer_time <= i_aer_time;
                    latched_aer_addr <= i_aer_addr;
                end

                S_COMPUTE: begin
                    // ִ��: t_i * W[i, j]
                    mult_result <= $signed(latched_aer_time) * $signed(i_bram_data);
                end
                
                S_SEND_DONE: begin
                    if (!i_reset_potential) begin // ���⸴λʱ���
                        V_j_reg <= V_j_reg + mult_result;
                    end
                end
            endcase
        end
    end

endmodule