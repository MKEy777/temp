`timescale 1ns / 1ps

/*
 * ģ��: SNN_Array_4PE [�ع���]
 * ����: 4-PE ��������
 * ְ��:
 * 1. ���� 4 x PE_GALS_Wrapper (ʹ�� CE)��
 * 2. ���� 1 x GALS_Collector_Unit��
 * 3. ʵ�� 32-bit -> 4x 8-bit Ȩ�ؽ������
 * 4. [���Ƴ�] BRAM ��ַƫ������ӡ�
 */
module SNN_Array_4PE #(
    parameter TIME_W   = 8,
    parameter WEIGHT_W = 8,
    parameter ADDR_W   = 10, // SNN ����ά��(160) + ƫ����
    parameter ACC_W    = 32
)(
    input  wire                 local_clk,
    input  wire                 rst_n,
    input  wire                 i_clk_en, // ** ����: ���м�ʱ��ʹ�� **

    // GALS �¼����� (�㲥)
    input  wire                 i_aer_req,
    input  wire signed [TIME_W-1:0] i_aer_time,
    input  wire [ADDR_W-1:0]        i_aer_addr,
    
    // SNN FSM ���Ʋ���
    // [���Ƴ�] i_bram_addr_offset
    input  wire signed [TIME_W-1:0] i_t_min,
    input  wire [3:0]               i_pe_enable,       // (PE ��ʱ��ʹ��)
    input  wire [3:0]               i_reset_potential,
    
    // ר�� BRAM �ӿ� (32-bit ��)
    output wire                 o_bram_en,
    // [���Ƴ�] o_bram_addr
    input  wire signed [31:0]   i_bram_data_32b,

    // GALS ���� (-> SNN_Engine)
    output wire                 o_array_aer_ack,
    output wire                 o_array_error, // (��¶ Collector ״̬)
    output wire                 o_array_busy,  // (��¶ Collector ״̬)

    // ��λ��� (-> SNN_Engine)
    output wire signed [4*ACC_W-1:0] o_potential_flat
);

    // �ڲ�����
    wire [3:0] pe_done_reqs;
    wire [3:0] pe_done_acks;
    wire [3:0] pe_bram_en_vec; // (���� 4 �� PE �� en �ź�)

    // ** �ؼ�: 32-bit -> 4x 8-bit Ȩ�ؽ���� **
    wire signed [WEIGHT_W-1:0] pe_weights [0:3]; 
    assign pe_weights[0] = i_bram_data_32b[ 7: 0]; // PE0 (LSB)
    assign pe_weights[1] = i_bram_data_32b[15: 8]; // PE1
    assign pe_weights[2] = i_bram_data_32b[23:16]; // PE2
    assign pe_weights[3] = i_bram_data_32b[31:24]; // PE3 (MSB)
    
    // --- 1. ���� 4-PE ���� (ʹ���ع���� PE) ---
    genvar i;
    generate
        for (i = 0; i < 4; i = i + 1) begin : gen_pe_array
            
            // ** ʵ�����ع���� PE (�� i_clk_en) **
            PE_GALS_Wrapper #(
                .TIME_W   ( TIME_W   ),
                .WEIGHT_W ( WEIGHT_W ),
                .ADDR_W   ( ADDR_W   ),
                .ACC_W    ( ACC_W    )
            ) pe_inst (
                .local_clk ( local_clk ),
                .rst_n     ( rst_n ),
                
                // ** �ؼ�: ������Ϻ��ʱ��ʹ�� **
                .i_clk_en  ( i_clk_en & i_pe_enable[i] ),
                
                .i_aer_req   ( i_aer_req ),
                .i_aer_time  ( i_aer_time ),
                .i_aer_addr  ( i_aer_addr ), // ��ֱַ��͸��
                .i_t_min     ( i_t_min ),
                
                .o_done_req ( pe_done_reqs[i] ),
                .i_done_ack ( pe_done_acks[i] ),
                
                .o_bram_en   ( pe_bram_en_vec[i] ),
                .i_bram_data ( pe_weights[i] ), // ���ӽ����� 8-bit Ȩ��
                
                .i_reset_potential ( i_reset_potential[i] ),
                .o_potential_j     ( o_potential_flat[(i+1)*ACC_W-1 -: ACC_W] )
            );
        end
    endgenerate

    // --- ���� BRAM ���� ---
    
    // [���Ƴ�] ��ַ���� (�� SNN_Engine ����)
    // assign o_bram_addr = i_aer_addr + i_bram_addr_offset; 
    
    // �κ�һ�����PE�����Դ���BRAM��ȡ
    assign o_bram_en = pe_bram_en_vec[0] | pe_bram_en_vec[1] |
                       pe_bram_en_vec[2] | pe_bram_en_vec[3];

    // --- 2. ���� GALS Collector (ʹ�����ṩ�İ汾) ---
    GALS_Collector_Unit #(
        .OUT_NEURONS ( 4 ),
        .WATCHDOG_TIMEOUT ( 10000 )
    ) collector_inst (
        .local_clk ( local_clk ),
        .rst_n     ( rst_n ),
        
        .i_aer_req ( i_aer_req ),
        .o_aer_ack ( o_array_aer_ack ),
        
        .i_pe_done_req_vec ( pe_done_reqs ),
        .o_pe_done_ack_vec ( pe_done_acks ),
        .o_error ( o_array_error ),
        .o_busy  ( o_array_busy )
    );

endmodule