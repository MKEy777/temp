`timescale 1ns / 1ps

/*
 * ģ��: ArgMax_Unit
 * ����: �ҳ� N ����λ�е����ֵ������
 * ����:
 * 1. VEC_LEN = 3 (���� train.py)
 * 2. DATA_W = 32 (ƥ�� PE_GALS_Wrapper �� 32-bit �ۼ���)
 */
module ArgMax_Unit #(
    parameter VEC_LEN = 3,  // ����� (���� train.py)
    parameter DATA_W  = 32  // �ؼ�: 32-bit (ƥ�� PE �ۼ���) 
) (
    input wire                        clk,
    input wire                        rst_n,
    input wire                        i_valid, // ���� SNN_Engine
    input wire signed [VEC_LEN*DATA_W-1:0] i_potentials_flat,

    output reg                        o_valid,
    output reg [$clog2(VEC_LEN)-1:0]  o_predicted_class
);

    // �ڲ��Ĵ��������ڱ��浱ǰ���ֵ�������� (����߼�)
    reg signed [DATA_W-1:0]     max_val;
    reg [$clog2(VEC_LEN)-1:0] max_idx;
    
    integer i;
    wire signed [DATA_W-1:0] potentials [0:VEC_LEN-1];

    // ��������λ
    genvar j;
    generate
        for (j = 0; j < VEC_LEN; j = j + 1) begin : unpack_potentials
            assign potentials[j] = i_potentials_flat[(j+1)*DATA_W-1 -: DATA_W];
        end
    endgenerate

    // ����߼�: Ѱ�����ֵ
    always @(*) begin
        max_val = potentials[0];
        max_idx = 0;
        
        for (i = 1; i < VEC_LEN; i = i + 1) begin
            if (potentials[i] > max_val) begin
                max_val = potentials[i];
                max_idx = i;
            end
        end
    end

    // ʱ���߼�: �Ĵ���
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            o_valid <= 1'b0;
            o_predicted_class <= 0;
        end else begin
            o_valid <= i_valid;
            if (i_valid) begin
                o_predicted_class <= max_idx;
            end
        end
    end

endmodule